module alphaDataMux(
	input [3:0] row,
	input [5:0] index,
	output wire [7:0] chardata
);

reg [4:0] data;

always @(row, index) begin
	case ({index,row})
		//@ 0
		10'b0000000010: data = 5'b01110;
		10'b0000000011: data = 5'b10001;
		10'b0000000100: data = 5'b00001;
		10'b0000000101: data = 5'b01101;
		10'b0000000110: data = 5'b10101;
		10'b0000000111: data = 5'b10101;
		10'b0000001000: data = 5'b01110;
		//A 1
		10'b0000010010: data = 5'b00100;
		10'b0000010011: data = 5'b01010;
		10'b0000010100: data = 5'b10001;
		10'b0000010101: data = 5'b10001;
		10'b0000010110: data = 5'b11111;
		10'b0000010111: data = 5'b10001;
		10'b0000011000: data = 5'b10000;
		//B 2
		10'b0000100010: data = 5'b11110;
		10'b0000100011: data = 5'b01001;
		10'b0000100100: data = 5'b01001;
		10'b0000100101: data = 5'b01110;
		10'b0000100110: data = 5'b01001;
		10'b0000100111: data = 5'b01001;
		10'b0000101000: data = 5'b11110;
		//C 3
		10'b0000110010: data = 5'b01110;
		10'b0000110011: data = 5'b10001;
		10'b0000110100: data = 5'b10000;
		10'b0000110101: data = 5'b10000;
		10'b0000110110: data = 5'b10000;
		10'b0000110111: data = 5'b10001;
		10'b0000111000: data = 5'b01110;
		//D 4
		10'b0001000010: data = 5'b11110;
		10'b0001000011: data = 5'b01001;
		10'b0001000100: data = 5'b01001;
		10'b0001000101: data = 5'b01001;
		10'b0001000110: data = 5'b01001;
		10'b0001000111: data = 5'b01001;
		10'b0001001000: data = 5'b11110;
		//E 5
		10'b0001010010: data = 5'b11111;
		10'b0001010011: data = 5'b10000;
		10'b0001010100: data = 5'b10000;
		10'b0001010101: data = 5'b11110;
		10'b0001010110: data = 5'b10000;
		10'b0001010111: data = 5'b10000;
		10'b0001011000: data = 5'b11111;
		//F 6
		10'b0001100010: data = 5'b11111;
		10'b0001100011: data = 5'b10000;
		10'b00011100100: data = 5'b10000;
		10'b0001100101: data = 5'b11110;
		10'b0001100110: data = 5'b10000;
		10'b00010100111: data = 5'b10000;
		10'b0001101000: data = 5'b10000;
		//G 7
		10'b0001110010: data = 5'b01111;
		10'b0001110011: data = 5'b10000;
		10'b0001110100: data = 5'b10000;
		10'b0001110101: data = 5'b10011;
		10'b0001110110: data = 5'b10001;
		10'b0001110111: data = 5'b10001;
		10'b0001111000: data = 5'b01110;
		//H 8
		10'b0010000010: data = 5'b10001;
		10'b0010000011: data = 5'b10001;
		10'b0010000100: data = 5'b10001;
		10'b0010000101: data = 5'b11111;
		10'b0010000110: data = 5'b10001;
		10'b0010000111: data = 5'b10001;
		10'b0010001000: data = 5'b10001;
		//I 9
		10'b0010010010: data = 5'b01110;
		10'b0010010011: data = 5'b00100;
		10'b0010010100: data = 5'b00100;
		10'b0010010101: data = 5'b00100;
		10'b0010010110: data = 5'b00100;
		10'b0010010111: data = 5'b00100;
		10'b0010011000: data = 5'b01110;
		//J 10
		10'b0010100010: data = 5'b00001;
		10'b0010100011: data = 5'b00001;
		10'b0010100100: data = 5'b00001;
		10'b0010100101: data = 5'b00001;
		10'b0010100110: data = 5'b10001;
		10'b0010100111: data = 5'b10001;
		10'b0010101000: data = 5'b01110;
		//K 11
		10'b0010110010: data = 5'b10001;
		10'b0010110011: data = 5'b10010;
		10'b0010110100: data = 5'b10100;
		10'b0010110101: data = 5'b11000;
		10'b0010110110: data = 5'b10100;
		10'b0010110111: data = 5'b10010;
		10'b0010111000: data = 5'b10001;
		//L 12
		10'b0011000010: data = 5'b10000;
		10'b0011000011: data = 5'b10000;
		10'b0011000100: data = 5'b10000;
		10'b0011000101: data = 5'b10000;
		10'b0011000110: data = 5'b10000;
		10'b0011000111: data = 5'b10000;
		10'b0011001000: data = 5'b11111;
		//M 13
		10'b0011010010: data = 5'b10001;
		10'b0011010011: data = 5'b11011;
		10'b0011010100: data = 5'b10101;
		10'b0011010101: data = 5'b10101;
		10'b0011010110: data = 5'b10001;
		10'b0011010111: data = 5'b10001;
		10'b0011011000: data = 5'b10001;
		//N 14
		10'b0011100010: data = 5'b10001;
		10'b0011100011: data = 5'b11001;
		10'b0011100100: data = 5'b10101;
		10'b0011100101: data = 5'b10011;
		10'b0011100110: data = 5'b10001;
		10'b0011100111: data = 5'b10001;
		10'b0011101000: data = 5'b10001;
		//O 15
		10'b0011110010: data = 5'b01110;
		10'b0011110011: data = 5'b10001;
		10'b0011110100: data = 5'b10001;
		10'b0011110101: data = 5'b10001;
		10'b0011110110: data = 5'b10001;
		10'b0011110111: data = 5'b10001;
		10'b0011111000: data = 5'b01110;
		//P 16
		10'b0100000010: data = 5'b11110;
		10'b0100000011: data = 5'b10001;
		10'b0100000100: data = 5'b10001;
		10'b0100000101: data = 5'b11110;
		10'b0100000110: data = 5'b10000;
		10'b0100000111: data = 5'b10000;
		10'b0100001000: data = 5'b10000;
		//Q 17
		10'b0100010010: data = 5'b01110;
		10'b0100010011: data = 5'b10001;
		10'b0100010100: data = 5'b10001;
		10'b0100010101: data = 5'b10001;
		10'b0100010110: data = 5'b10101;
		10'b0100010111: data = 5'b10010;
		10'b0100011000: data = 5'b01101;
		//R 18
		10'b0100100010: data = 5'b11110;
		10'b0100100011: data = 5'b10001;
		10'b0100100100: data = 5'b10001;
		10'b0100100101: data = 5'b11110;
		10'b0100100110: data = 5'b10100;
		10'b0100100111: data = 5'b10010;
		10'b0100101000: data = 5'b10001;
		//S 19
		10'b0100110010: data = 5'b01110;
		10'b0100110011: data = 5'b10001;
		10'b0100110100: data = 5'b01000;
		10'b0100110101: data = 5'b00100;
		10'b0100110110: data = 5'b00010;
		10'b0100110111: data = 5'b10001;
		10'b0100111000: data = 5'b01110;
		//T 20
		10'b0101000010: data = 5'b11111;
		10'b0101000011: data = 5'b00100;
		10'b0101000100: data = 5'b00100;
		10'b0101000101: data = 5'b00100;
		10'b0101000110: data = 5'b00100;
		10'b0101000111: data = 5'b00100;
		10'b0101001000: data = 5'b00100;
		//U 21
		10'b0101010010: data = 5'b10001;
		10'b0101010011: data = 5'b10001;
		10'b0101010100: data = 5'b10001;
		10'b0101010101: data = 5'b10001;
		10'b0101010110: data = 5'b10001;
		10'b0101010111: data = 5'b10001;
		10'b0101011000: data = 5'b01110;
		//V 22
		10'b0101100010: data = 5'b10001;
		10'b0101100011: data = 5'b10001;
		10'b0101100100: data = 5'b10001;
		10'b0101100101: data = 5'b01010;
		10'b0101100110: data = 5'b01010;
		10'b0101100111: data = 5'b00100;
		10'b0101101000: data = 5'b00100;
		//W 23
		10'b0101110010: data = 5'b10001;
		10'b0101110011: data = 5'b10001;
		10'b0101110100: data = 5'b10001;
		10'b0101110101: data = 5'b10101;
		10'b0101110110: data = 5'b10101;
		10'b0101110111: data = 5'b11011;
		10'b0101111000: data = 5'b10001;
		//X 24
		10'b0110000010: data = 5'b10001;
		10'b0110000011: data = 5'b10001;
		10'b0110000100: data = 5'b01010;
		10'b0110000101: data = 5'b00100;
		10'b0110000110: data = 5'b01010;
		10'b0110000111: data = 5'b10001;
		10'b0110001000: data = 5'b10001;
		//Y 25
		10'b0110010010: data = 5'b10001;
		10'b0110010011: data = 5'b10001;
		10'b0110010100: data = 5'b01010;
		10'b0110010101: data = 5'b00100;
		10'b0110010110: data = 5'b00100;
		10'b0110010111: data = 5'b00100;
		10'b0110011000: data = 5'b00100;
		//Z 26
		10'b0110100010: data = 5'b11111;
		10'b0110100011: data = 5'b00001;
		10'b0110100100: data = 5'b00010;
		10'b0110100101: data = 5'b00100;
		10'b0110100110: data = 5'b01000;
		10'b0110100111: data = 5'b10000;
		10'b0110101000: data = 5'b11111;
		//[ 27
		10'b0110110010: data = 5'b11100;
		10'b0110110011: data = 5'b10000;
		10'b0110110100: data = 5'b10000;
		10'b0110110101: data = 5'b10000;
		10'b0110110110: data = 5'b10000;
		10'b0110110111: data = 5'b10000;
		10'b0110111000: data = 5'b11100;
		// \ 28
		10'b0111000010: data = 5'b11100;
		10'b0111000011: data = 5'b10000;
		10'b0111000100: data = 5'b10000;
		10'b0111000101: data = 5'b10000;
		10'b0111000110: data = 5'b10000;
		10'b0111000111: data = 5'b10000;
		10'b0111001000: data = 5'b11100;
		// ] 29
		10'b0111010010: data = 5'b11100;
		10'b0111010011: data = 5'b10000;
		10'b0111010100: data = 5'b10000;
		10'b0111010101: data = 5'b10000;
		10'b0111010110: data = 5'b10000;
		10'b0111010111: data = 5'b10000;
		10'b0111011000: data = 5'b11100;
		// (up) 30
		10'b0111100010: data = 5'b00100;
		10'b0111100011: data = 5'b01110;
		10'b0111100100: data = 5'b10101;
		10'b0111100101: data = 5'b00100;
		10'b0111100110: data = 5'b00100;
		10'b0111100111: data = 5'b00100;
		10'b0111101000: data = 5'b00100;
		// (left) 31
		10'b0111110010: data = 5'b00000;
		10'b0111110011: data = 5'b00100;
		10'b0111110100: data = 5'b01000;
		10'b0111110101: data = 5'b11111;
		10'b0111110110: data = 5'b01000;
		10'b0111110111: data = 5'b00100;
		10'b0111111000: data = 5'b00000;
		// (space) 32
		10'b1000000010: data = 5'b00000;
		10'b1000000011: data = 5'b00000;
		10'b1000000100: data = 5'b00000;
		10'b1000000101: data = 5'b00000;
		10'b1000000110: data = 5'b00000;
		10'b1000000111: data = 5'b00000;
		10'b1000001000: data = 5'b00000;
		// ! 33
		10'b1000010010: data = 5'b00100;
		10'b1000010011: data = 5'b00100;
		10'b1000010100: data = 5'b00100;
		10'b1000010101: data = 5'b00100;
		10'b1000010110: data = 5'b00100;
		10'b1000010111: data = 5'b00000;
		10'b1000011000: data = 5'b00100;
		// " 34
		10'b1000100010: data = 5'b01010;
		10'b1000100011: data = 5'b01010;
		10'b1000100100: data = 5'b00000;
		10'b1000100101: data = 5'b00000;
		10'b1000100110: data = 5'b00000;
		10'b1000100111: data = 5'b00000;
		10'b1000101000: data = 5'b00000;
		// # 35
		10'b1000110010: data = 5'b01010;
		10'b1000110011: data = 5'b01010;
		10'b1000110100: data = 5'b11011;
		10'b1000110101: data = 5'b00000;
		10'b1000110110: data = 5'b11011;
		10'b1000110111: data = 5'b01010;
		10'b1000111000: data = 5'b01010;
		// $ 36
		10'b1001000010: data = 5'b00100;
		10'b1001000011: data = 5'b01111;
		10'b1001000100: data = 5'b10000;
		10'b1001000101: data = 5'b01110;
		10'b1001000110: data = 5'b00001;
		10'b1001000111: data = 5'b11110;
		10'b1001001000: data = 5'b00100;
		// % 37
		10'b1001010010: data = 5'b11001;
		10'b1001010011: data = 5'b11001;
		10'b1001010100: data = 5'b00010;
		10'b1001010101: data = 5'b00100;
		10'b1001010110: data = 5'b01000;
		10'b1001010111: data = 5'b10011;
		10'b1001011000: data = 5'b10011;
		// & 38
		10'b1001100010: data = 5'b01000;
		10'b1001100011: data = 5'b10100;
		10'b1001100100: data = 5'b10100;
		10'b1001100101: data = 5'b01000;
		10'b1001100110: data = 5'b10101;
		10'b1001100111: data = 5'b10010;
		10'b1001101000: data = 5'b01101;
		// ' 39
		10'b1001110010: data = 5'b01100;
		10'b1001110011: data = 5'b01100;
		10'b1001110100: data = 5'b01100;
		10'b1001110101: data = 5'b00000;
		10'b1001110110: data = 5'b00000;
		10'b1001110111: data = 5'b00000;
		10'b1001111000: data = 5'b00000;
		// ( 40
		10'b1010000010: data = 5'b00100;
		10'b1010000011: data = 5'b01000;
		10'b1010000100: data = 5'b10000;
		10'b1010000101: data = 5'b10000;
		10'b1010000110: data = 5'b10000;
		10'b1010000111: data = 5'b01000;
		10'b1010001000: data = 5'b00100;
		// ) 41
		10'b1010010010: data = 5'b00100;
		10'b1010010011: data = 5'b00010;
		10'b1010010100: data = 5'b00001;
		10'b1010010101: data = 5'b00001;
		10'b1010010110: data = 5'b00001;
		10'b1010010111: data = 5'b00010;
		10'b1010011000: data = 5'b00100;
		// * 42
		10'b1010100010: data = 5'b00000;
		10'b1010100011: data = 5'b00100;
		10'b1010100100: data = 5'b01110;
		10'b1010100101: data = 5'b11111;
		10'b1010100110: data = 5'b01110;
		10'b1010100111: data = 5'b00100;
		10'b1010101000: data = 5'b00000;
		// + 43
		10'b1010110010: data = 5'b00000;
		10'b1010110011: data = 5'b00100;
		10'b1010110100: data = 5'b00100;
		10'b1010110101: data = 5'b11111;
		10'b1010110110: data = 5'b00100;
		10'b1010110111: data = 5'b00100;
		10'b1010111000: data = 5'b00000;
		// , 44
		10'b1011000010: data = 5'b00000;
		10'b1011000011: data = 5'b00000;
		10'b1011000100: data = 5'b00000;
		10'b1011000101: data = 5'b11000;
		10'b1011000110: data = 5'b11000;
		10'b1011000111: data = 5'b01000;
		10'b1011001000: data = 5'b10000;
		// - 45
		10'b1011010010: data = 5'b00000;
		10'b1011010011: data = 5'b00000;
		10'b1011010100: data = 5'b00000;
		10'b1011010101: data = 5'b11111;
		10'b1011010110: data = 5'b00000;
		10'b1011010111: data = 5'b00000;
		10'b1011011000: data = 5'b00000;
		// . 46
		10'b1011100010: data = 5'b00000;
		10'b1011100011: data = 5'b00000;
		10'b1011100100: data = 5'b00000;
		10'b1011100101: data = 5'b00000;
		10'b1011100110: data = 5'b00000;
		10'b1011100111: data = 5'b11000;
		10'b1011101000: data = 5'b11000;
		// / 47
		10'b1011110010: data = 5'b00001;
		10'b1011110011: data = 5'b00001;
		10'b1011110100: data = 5'b00010;
		10'b1011110101: data = 5'b00100;
		10'b1011110110: data = 5'b01000;
		10'b1011110111: data = 5'b10000;
		10'b1011111000: data = 5'b10000;
		// 0 48
		10'b1100000010: data = 5'b01100;
		10'b1100000011: data = 5'b10010;
		10'b1100000100: data = 5'b10010;
		10'b1100000101: data = 5'b10010;
		10'b1100000110: data = 5'b10010;
		10'b1100000111: data = 5'b10010;
		10'b1100001000: data = 5'b01100;
		// 1 49
		10'b1100010010: data = 5'b00100;
		10'b1100010011: data = 5'b01100;
		10'b1100010100: data = 5'b00100;
		10'b1100010101: data = 5'b00100;
		10'b1100010110: data = 5'b00100;
		10'b1100010111: data = 5'b00100;
		10'b1100011000: data = 5'b01110;
		// 2 50
		10'b1100100010: data = 5'b01110;
		10'b1100100011: data = 5'b10001;
		10'b1100100100: data = 5'b00001;
		10'b1100100101: data = 5'b01110;
		10'b1100100110: data = 5'b10000;
		10'b1100100111: data = 5'b10000;
		10'b1100101000: data = 5'b11111;
		// 3 51
		10'b1100110010: data = 5'b01110;
		10'b1100110011: data = 5'b10001;
		10'b1100110100: data = 5'b00001;
		10'b1100110101: data = 5'b00110;
		10'b1100110110: data = 5'b00001;
		10'b1100110111: data = 5'b10001;
		10'b1100111000: data = 5'b01110;
		// 4 52
		10'b1101000010: data = 5'b00010;
		10'b1101000011: data = 5'b00110;
		10'b1101000100: data = 5'b01010;
		10'b1101000101: data = 5'b11110;
		10'b1101000110: data = 5'b00010;
		10'b1101000111: data = 5'b00010;
		10'b1101001000: data = 5'b00010;
		// 5 53
		10'b1101010010: data = 5'b11111;
		10'b1101010011: data = 5'b10000;
		10'b1101010100: data = 5'b10000;
		10'b1101010101: data = 5'b11110;
		10'b1101010110: data = 5'b00001;
		10'b1101010111: data = 5'b10001;
		10'b1101011000: data = 5'b01110;
		// 6 54
		10'b1101100010: data = 5'b01110;
		10'b1101100011: data = 5'b10000;
		10'b1101100100: data = 5'b10000;
		10'b1101100101: data = 5'b11110;
		10'b1101100110: data = 5'b10001;
		10'b1101100111: data = 5'b10001;
		10'b1101101000: data = 5'b01110;
		// 7 55
		10'b1101110010: data = 5'b11111;
		10'b1101110011: data = 5'b00001;
		10'b1101110100: data = 5'b00010;
		10'b1101110101: data = 5'b00100;
		10'b1101110110: data = 5'b01000;
		10'b1101110111: data = 5'b10000;
		10'b1101111000: data = 5'b10000;
		// 8 56
		10'b1110000010: data = 5'b01110;
		10'b1110000011: data = 5'b10001;
		10'b1110000100: data = 5'b10001;
		10'b1110000101: data = 5'b01110;
		10'b1110000110: data = 5'b10001;
		10'b1110000111: data = 5'b10001;
		10'b1110001000: data = 5'b01110;
		// 9 57
		10'b1110010010: data = 5'b01110;
		10'b1110010011: data = 5'b10001;
		10'b1110010100: data = 5'b10001;
		10'b1110010101: data = 5'b01111;
		10'b1110010110: data = 5'b00001;
		10'b1110010111: data = 5'b00001;
		10'b1110011000: data = 5'b01110;
		// : 58
		10'b1110100010: data = 5'b00000;
		10'b1110100011: data = 5'b01100;
		10'b1110100100: data = 5'b01100;
		10'b1110100101: data = 5'b00000;
		10'b1110100110: data = 5'b01100;
		10'b1110100111: data = 5'b01100;
		10'b1110101000: data = 5'b00000;
		// ; 59
		10'b1110110010: data = 5'b01100;
		10'b1110110011: data = 5'b01100;
		10'b1110110100: data = 5'b00000;
		10'b1110110101: data = 5'b01100;
		10'b1110110110: data = 5'b01100;
		10'b1110110111: data = 5'b00100;
		10'b1110111000: data = 5'b01000;
		// < 60
		10'b1111000010: data = 5'b00010;
		10'b1111000011: data = 5'b00100;
		10'b1111000100: data = 5'b01000;
		10'b1111000101: data = 5'b10000;
		10'b1111000110: data = 5'b01000;
		10'b1111000111: data = 5'b00100;
		10'b1111001000: data = 5'b00010;
		// = 61
		10'b1111010010: data = 5'b00000;
		10'b1111010011: data = 5'b00000;
		10'b1111010100: data = 5'b11111;
		10'b1111010101: data = 5'b10000;
		10'b1111010110: data = 5'b11111;
		10'b1111010111: data = 5'b00000;
		10'b1111011000: data = 5'b00010;
		// > 62
		10'b1111100010: data = 5'b01000;
		10'b1111100011: data = 5'b00100;
		10'b1111100100: data = 5'b00010;
		10'b1111100101: data = 5'b00001;
		10'b1111100110: data = 5'b00010;
		10'b1111100111: data = 5'b00100;
		10'b1111101000: data = 5'b01000;
		// ? 63
		10'b1111110010: data = 5'b01100;
		10'b1111110011: data = 5'b10010;
		10'b1111110100: data = 5'b00010;
		10'b1111110101: data = 5'b00100;
		10'b1111110110: data = 5'b00100;
		10'b1111110111: data = 5'b00000;
		10'b1111111000: data = 5'b00100;
		// 
		default: data = 5'd0;
	endcase
end

assign chardata = {2'b00,data,1'b0};

endmodule
/*
Tested working in simulation
*/